
module part3 ( clk, reset, a, valid_in, g, valid_out );
  input [7:0] a;
  output [9:0] g;
  input clk, reset, valid_in;
  output valid_out;
  wire   enable_f, enable_g, N3, N4, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n59, n60, n63, n64, n65, n66, n68, n69, n70, n71,
         n72, n73, n74, n76, n77, n80, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685;
  wire   [7:0] a_reg;
  wire   [19:0] f;

  DFF_X1 \f_reg[0]  ( .D(n55), .CK(clk), .Q(f[0]), .QN(n668) );
  DFF_X1 enable_f_reg ( .D(N3), .CK(clk), .Q(enable_f), .QN(n666) );
  DFF_X1 \f_reg[1]  ( .D(n56), .CK(clk), .Q(f[1]), .QN(n664) );
  DFF_X1 \a_reg_reg[7]  ( .D(n680), .CK(clk), .Q(n660), .QN(a_reg[7]) );
  DFF_X1 \a_reg_reg[6]  ( .D(n681), .CK(clk), .Q(n659), .QN(a_reg[6]) );
  DFF_X1 \a_reg_reg[4]  ( .D(n682), .CK(clk), .Q(n661), .QN(a_reg[4]) );
  DFF_X1 \a_reg_reg[3]  ( .D(n683), .CK(clk), .Q(n662), .QN(a_reg[3]) );
  DFF_X1 \a_reg_reg[0]  ( .D(n684), .CK(clk), .Q(n667), .QN(a_reg[0]) );
  DFF_X1 \f_reg[2]  ( .D(n679), .CK(clk), .Q(n651), .QN(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(n678), .CK(clk), .Q(n669), .QN(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(n59), .CK(clk), .Q(f[4]), .QN(n652) );
  DFF_X1 \f_reg[5]  ( .D(n60), .CK(clk), .Q(f[5]), .QN(n663) );
  DFF_X1 \f_reg[6]  ( .D(n677), .CK(clk), .Q(n653), .QN(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(n676), .CK(clk), .Q(n665), .QN(f[7]) );
  DFF_X1 \f_reg[8]  ( .D(n63), .CK(clk), .Q(f[8]), .QN(n654) );
  DFF_X1 \f_reg[10]  ( .D(n65), .CK(clk), .Q(f[10]), .QN(n650) );
  DFF_X1 \f_reg[12]  ( .D(n675), .CK(clk), .Q(n657), .QN(f[12]) );
  DFF_X1 \f_reg[13]  ( .D(n68), .CK(clk), .Q(f[13]), .QN(n670) );
  DFF_X1 \f_reg[14]  ( .D(n69), .CK(clk), .Q(f[14]), .QN(n658) );
  DFF_X1 \f_reg[15]  ( .D(n70), .CK(clk), .Q(f[15]), .QN(n648) );
  DFF_X1 \f_reg[16]  ( .D(n71), .CK(clk), .Q(f[16]), .QN(n656) );
  DFF_X1 \f_reg[17]  ( .D(n72), .CK(clk), .Q(f[17]), .QN(n671) );
  DFF_X1 \f_reg[18]  ( .D(n73), .CK(clk), .Q(f[18]), .QN(n655) );
  DFF_X1 \f_reg[19]  ( .D(n74), .CK(clk), .Q(f[19]), .QN(n649) );
  DFF_X1 enable_out_reg ( .D(n685), .CK(clk), .Q(valid_out) );
  DFF_X1 enable_g_reg ( .D(N4), .CK(clk), .Q(enable_g) );
  DFF_X1 \g_reg[9]  ( .D(n54), .CK(clk), .Q(g[9]) );
  DFF_X1 \a_reg_reg[2]  ( .D(n77), .CK(clk), .Q(a_reg[2]), .QN(n674) );
  DFF_X1 \a_reg_reg[1]  ( .D(n76), .CK(clk), .Q(a_reg[1]), .QN(n673) );
  DFF_X1 \a_reg_reg[5]  ( .D(n80), .CK(clk), .Q(a_reg[5]), .QN(n672) );
  DFF_X1 \g_reg[8]  ( .D(n53), .CK(clk), .Q(g[8]) );
  DFF_X1 \g_reg[7]  ( .D(n52), .CK(clk), .Q(g[7]) );
  DFF_X1 \f_reg[9]  ( .D(n64), .CK(clk), .Q(f[9]) );
  DFF_X1 \g_reg[6]  ( .D(n51), .CK(clk), .Q(g[6]) );
  DFF_X1 \f_reg[11]  ( .D(n66), .CK(clk), .Q(f[11]) );
  DFF_X1 \g_reg[5]  ( .D(n50), .CK(clk), .Q(g[5]) );
  DFF_X1 \g_reg[4]  ( .D(n49), .CK(clk), .Q(g[4]) );
  DFF_X1 \g_reg[3]  ( .D(n48), .CK(clk), .Q(g[3]) );
  DFF_X1 \g_reg[2]  ( .D(n47), .CK(clk), .Q(g[2]) );
  DFF_X1 \g_reg[1]  ( .D(n46), .CK(clk), .Q(g[1]) );
  DFF_X1 \g_reg[0]  ( .D(n45), .CK(clk), .Q(g[0]) );
  INV_X1 U88 ( .A(n300), .ZN(n577) );
  INV_X1 U89 ( .A(n475), .ZN(n527) );
  INV_X1 U90 ( .A(n393), .ZN(n529) );
  AOI21_X2 U91 ( .B1(n373), .B2(n83), .A(n338), .ZN(n574) );
  NAND2_X1 U92 ( .A1(n103), .A2(n102), .ZN(n326) );
  INV_X1 U93 ( .A(N4), .ZN(n294) );
  NOR2_X2 U94 ( .A1(f[18]), .A2(f[19]), .ZN(n616) );
  INV_X1 U95 ( .A(n254), .ZN(n307) );
  XNOR2_X1 U96 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U97 ( .A1(n484), .A2(n483), .ZN(n485) );
  AOI21_X1 U98 ( .B1(n503), .B2(n482), .A(n481), .ZN(n486) );
  NOR2_X1 U99 ( .A1(n378), .A2(n616), .ZN(n375) );
  NOR2_X1 U100 ( .A1(n322), .A2(n321), .ZN(n323) );
  XNOR2_X1 U101 ( .A(n539), .B(n538), .ZN(n541) );
  NOR2_X1 U102 ( .A1(n476), .A2(n537), .ZN(n538) );
  OAI21_X1 U103 ( .B1(n598), .B2(n543), .A(n544), .ZN(n539) );
  XNOR2_X1 U104 ( .A(n478), .B(n477), .ZN(n480) );
  INV_X1 U105 ( .A(n503), .ZN(n477) );
  INV_X1 U106 ( .A(n514), .ZN(n612) );
  XNOR2_X1 U107 ( .A(n494), .B(n87), .ZN(n496) );
  NAND2_X1 U108 ( .A1(n394), .A2(n447), .ZN(n458) );
  NAND2_X1 U109 ( .A1(n448), .A2(n450), .ZN(n394) );
  NOR2_X1 U110 ( .A1(n495), .A2(n326), .ZN(n498) );
  NAND2_X1 U111 ( .A1(n432), .A2(n616), .ZN(n428) );
  OAI21_X1 U112 ( .B1(n475), .B2(n474), .A(n473), .ZN(n540) );
  INV_X1 U113 ( .A(n463), .ZN(n474) );
  NAND2_X1 U114 ( .A1(n475), .A2(n472), .ZN(n473) );
  XNOR2_X1 U115 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U116 ( .A(n346), .B(n345), .ZN(n348) );
  MUX2_X1 U117 ( .A(n364), .B(n363), .S(n574), .Z(n416) );
  NOR2_X1 U118 ( .A1(n360), .A2(n359), .ZN(n361) );
  XNOR2_X1 U119 ( .A(n554), .B(n553), .ZN(n556) );
  NAND2_X1 U120 ( .A1(n552), .A2(n551), .ZN(n553) );
  OAI21_X1 U121 ( .B1(n560), .B2(n557), .A(n549), .ZN(n554) );
  NOR2_X1 U122 ( .A1(n575), .A2(n574), .ZN(n563) );
  AOI22_X1 U123 ( .A1(n532), .A2(n531), .B1(n530), .B2(n529), .ZN(n533) );
  NOR2_X1 U124 ( .A1(n528), .A2(n475), .ZN(n531) );
  XNOR2_X1 U125 ( .A(n356), .B(n355), .ZN(n358) );
  NAND2_X1 U126 ( .A1(n354), .A2(n353), .ZN(n355) );
  OAI21_X1 U127 ( .B1(n362), .B2(n360), .A(n351), .ZN(n356) );
  OAI21_X1 U128 ( .B1(n456), .B2(n560), .A(n455), .ZN(n598) );
  OR2_X1 U129 ( .A1(n557), .A2(n453), .ZN(n456) );
  INV_X1 U130 ( .A(n552), .ZN(n453) );
  NAND2_X1 U131 ( .A1(n460), .A2(n574), .ZN(n464) );
  NOR2_X1 U132 ( .A1(n460), .A2(n574), .ZN(n465) );
  NAND2_X1 U133 ( .A1(n509), .A2(n616), .ZN(n505) );
  NOR2_X1 U134 ( .A1(n509), .A2(n616), .ZN(n504) );
  XNOR2_X1 U135 ( .A(n318), .B(n317), .ZN(n320) );
  NAND2_X1 U136 ( .A1(n316), .A2(n315), .ZN(n317) );
  OAI21_X1 U137 ( .B1(n329), .B2(n322), .A(n313), .ZN(n318) );
  NAND2_X1 U138 ( .A1(n366), .A2(n86), .ZN(n367) );
  INV_X1 U139 ( .A(n372), .ZN(n366) );
  NAND2_X1 U140 ( .A1(n341), .A2(n387), .ZN(n401) );
  NAND2_X1 U141 ( .A1(n388), .A2(n390), .ZN(n341) );
  AND2_X1 U142 ( .A1(n378), .A2(n616), .ZN(n374) );
  OAI21_X1 U143 ( .B1(n329), .B2(n328), .A(n327), .ZN(n332) );
  AND2_X1 U144 ( .A1(n368), .A2(n326), .ZN(n372) );
  OAI21_X1 U145 ( .B1(n362), .B2(n311), .A(n310), .ZN(n373) );
  OR2_X1 U146 ( .A1(n360), .A2(n309), .ZN(n311) );
  AOI21_X1 U147 ( .B1(n353), .B2(n359), .A(n352), .ZN(n310) );
  INV_X1 U148 ( .A(n257), .ZN(n569) );
  NAND2_X1 U149 ( .A1(n573), .A2(n90), .ZN(n581) );
  OAI21_X1 U150 ( .B1(n626), .B2(n619), .A(n618), .ZN(n628) );
  NAND2_X1 U151 ( .A1(n624), .A2(n326), .ZN(n619) );
  AOI21_X1 U152 ( .B1(n617), .B2(n616), .A(n615), .ZN(n618) );
  OAI21_X1 U153 ( .B1(n503), .B2(n89), .A(n502), .ZN(n508) );
  NOR2_X1 U154 ( .A1(n501), .A2(n500), .ZN(n502) );
  NOR2_X1 U155 ( .A1(f[16]), .A2(f[17]), .ZN(n129) );
  INV_X1 U156 ( .A(n458), .ZN(n466) );
  OR2_X1 U157 ( .A1(n524), .A2(n527), .ZN(n521) );
  INV_X1 U158 ( .A(n401), .ZN(n404) );
  INV_X1 U159 ( .A(n405), .ZN(n407) );
  INV_X1 U160 ( .A(n606), .ZN(n607) );
  NAND2_X1 U161 ( .A1(n462), .A2(n300), .ZN(n544) );
  AND2_X1 U162 ( .A1(n555), .A2(n574), .ZN(n550) );
  OR2_X1 U163 ( .A1(n555), .A2(n574), .ZN(n552) );
  NAND2_X1 U164 ( .A1(n487), .A2(n569), .ZN(n483) );
  OR2_X1 U165 ( .A1(n391), .A2(n574), .ZN(n388) );
  NAND2_X1 U166 ( .A1(n391), .A2(n574), .ZN(n387) );
  AND2_X1 U167 ( .A1(n301), .A2(n343), .ZN(n362) );
  NAND2_X1 U168 ( .A1(n344), .A2(n346), .ZN(n301) );
  AOI21_X1 U169 ( .B1(n257), .B2(n185), .A(n181), .ZN(n267) );
  AOI21_X1 U170 ( .B1(n257), .B2(n658), .A(n648), .ZN(n181) );
  XNOR2_X1 U171 ( .A(n592), .B(n591), .ZN(n594) );
  NAND2_X1 U172 ( .A1(n585), .A2(n584), .ZN(n592) );
  NAND2_X1 U173 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U174 ( .A(n487), .ZN(n412) );
  INV_X1 U175 ( .A(n375), .ZN(n336) );
  NAND2_X1 U176 ( .A1(n312), .A2(n316), .ZN(n328) );
  AND2_X1 U177 ( .A1(n255), .A2(n303), .ZN(n329) );
  AOI21_X1 U178 ( .B1(n321), .B2(n316), .A(n314), .ZN(n327) );
  NOR2_X1 U179 ( .A1(n333), .A2(n616), .ZN(n331) );
  AOI22_X1 U180 ( .A1(n580), .A2(n579), .B1(n578), .B2(n577), .ZN(n582) );
  AND2_X1 U181 ( .A1(n575), .A2(n574), .ZN(n580) );
  INV_X1 U182 ( .A(n576), .ZN(n579) );
  NAND2_X1 U183 ( .A1(n542), .A2(n257), .ZN(n573) );
  AND2_X1 U184 ( .A1(n570), .A2(n569), .ZN(n571) );
  AND2_X1 U185 ( .A1(n568), .A2(n567), .ZN(n572) );
  NOR2_X1 U186 ( .A1(n576), .A2(n563), .ZN(n564) );
  XNOR2_X1 U187 ( .A(n602), .B(n601), .ZN(n604) );
  NOR2_X1 U188 ( .A1(n600), .A2(n599), .ZN(n601) );
  AOI21_X1 U189 ( .B1(n598), .B2(n586), .A(n597), .ZN(n602) );
  NOR2_X1 U190 ( .A1(n617), .A2(n616), .ZN(n626) );
  NAND2_X1 U191 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U192 ( .A(n422), .B(n421), .ZN(n424) );
  NOR2_X1 U193 ( .A1(n613), .A2(n616), .ZN(n605) );
  AND2_X1 U194 ( .A1(n613), .A2(n616), .ZN(n606) );
  AOI21_X1 U195 ( .B1(n598), .B2(n493), .A(n492), .ZN(n609) );
  NOR2_X1 U196 ( .A1(n595), .A2(n491), .ZN(n493) );
  OAI21_X1 U197 ( .B1(n596), .B2(n491), .A(n490), .ZN(n492) );
  OR2_X1 U198 ( .A1(n599), .A2(n489), .ZN(n491) );
  AOI21_X1 U199 ( .B1(n396), .B2(n458), .A(n395), .ZN(n503) );
  OAI21_X1 U200 ( .B1(n464), .B2(n467), .A(n468), .ZN(n395) );
  INV_X1 U201 ( .A(n435), .ZN(n441) );
  OAI21_X1 U202 ( .B1(n438), .B2(n504), .A(n505), .ZN(n439) );
  INV_X1 U203 ( .A(n500), .ZN(n438) );
  NAND2_X1 U204 ( .A1(n413), .A2(n484), .ZN(n497) );
  OR2_X1 U205 ( .A1(n498), .A2(n504), .ZN(n435) );
  XNOR2_X1 U206 ( .A(n431), .B(n430), .ZN(n433) );
  NAND2_X1 U207 ( .A1(n429), .A2(n428), .ZN(n430) );
  INV_X1 U208 ( .A(n380), .ZN(n381) );
  XNOR2_X1 U209 ( .A(n377), .B(n376), .ZN(n379) );
  AOI21_X1 U210 ( .B1(n401), .B2(n350), .A(n349), .ZN(n427) );
  NOR2_X1 U211 ( .A1(n403), .A2(n405), .ZN(n350) );
  OAI21_X1 U212 ( .B1(n402), .B2(n405), .A(n406), .ZN(n349) );
  NAND2_X1 U213 ( .A1(n84), .A2(n365), .ZN(n426) );
  INV_X1 U214 ( .A(n419), .ZN(n365) );
  INV_X1 U215 ( .A(n331), .ZN(n269) );
  AND2_X1 U216 ( .A1(n333), .A2(n616), .ZN(n330) );
  NAND2_X1 U217 ( .A1(f[18]), .A2(n649), .ZN(n103) );
  OAI21_X1 U218 ( .B1(n466), .B2(n465), .A(n464), .ZN(n471) );
  NAND2_X1 U219 ( .A1(n469), .A2(n468), .ZN(n470) );
  OR2_X1 U220 ( .A1(n347), .A2(n577), .ZN(n344) );
  NAND2_X1 U221 ( .A1(n347), .A2(n577), .ZN(n343) );
  XNOR2_X1 U222 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U223 ( .A(n459), .B(n466), .ZN(n461) );
  NOR2_X1 U224 ( .A1(n457), .A2(n465), .ZN(n459) );
  INV_X1 U225 ( .A(n464), .ZN(n457) );
  XNOR2_X1 U226 ( .A(n523), .B(n522), .ZN(n525) );
  NAND2_X1 U227 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U228 ( .A1(n530), .A2(n529), .ZN(n528) );
  XNOR2_X1 U229 ( .A(n401), .B(n398), .ZN(n400) );
  NOR2_X1 U230 ( .A1(n588), .A2(n600), .ZN(n589) );
  XNOR2_X1 U231 ( .A(n306), .B(n305), .ZN(n308) );
  INV_X1 U232 ( .A(n359), .ZN(n351) );
  INV_X1 U233 ( .A(n352), .ZN(n354) );
  AND2_X1 U234 ( .A1(n593), .A2(n326), .ZN(n583) );
  OR2_X1 U235 ( .A1(n593), .A2(n326), .ZN(n584) );
  AND2_X1 U236 ( .A1(n547), .A2(n577), .ZN(n543) );
  AND2_X1 U237 ( .A1(n540), .A2(n567), .ZN(n537) );
  AND2_X1 U238 ( .A1(n561), .A2(n529), .ZN(n558) );
  NOR2_X1 U239 ( .A1(n561), .A2(n529), .ZN(n557) );
  AND2_X1 U240 ( .A1(n454), .A2(n520), .ZN(n560) );
  NAND2_X1 U241 ( .A1(n521), .A2(n523), .ZN(n454) );
  OR2_X1 U242 ( .A1(n451), .A2(n529), .ZN(n448) );
  NAND2_X1 U243 ( .A1(n451), .A2(n529), .ZN(n447) );
  XNOR2_X1 U244 ( .A(n390), .B(n389), .ZN(n392) );
  NAND2_X1 U245 ( .A1(n479), .A2(n567), .ZN(n482) );
  XNOR2_X1 U246 ( .A(n409), .B(n408), .ZN(n411) );
  NAND2_X1 U247 ( .A1(n407), .A2(n406), .ZN(n408) );
  OAI21_X1 U248 ( .B1(n404), .B2(n403), .A(n402), .ZN(n409) );
  NOR2_X1 U249 ( .A1(n414), .A2(n419), .ZN(n415) );
  INV_X1 U250 ( .A(n312), .ZN(n322) );
  INV_X1 U251 ( .A(n321), .ZN(n313) );
  INV_X1 U252 ( .A(n314), .ZN(n315) );
  AND2_X1 U253 ( .A1(n363), .A2(n567), .ZN(n359) );
  AND2_X1 U254 ( .A1(n357), .A2(n569), .ZN(n352) );
  NOR2_X1 U255 ( .A1(n357), .A2(n569), .ZN(n309) );
  NOR2_X1 U256 ( .A1(n363), .A2(n567), .ZN(n360) );
  INV_X1 U257 ( .A(n309), .ZN(n353) );
  OR2_X1 U258 ( .A1(n324), .A2(n569), .ZN(n312) );
  AND2_X1 U259 ( .A1(n324), .A2(n569), .ZN(n321) );
  AND2_X1 U260 ( .A1(n319), .A2(n326), .ZN(n314) );
  OR2_X1 U261 ( .A1(n319), .A2(n326), .ZN(n316) );
  INV_X1 U262 ( .A(n267), .ZN(n182) );
  NOR2_X1 U263 ( .A1(n578), .A2(n577), .ZN(n576) );
  OAI21_X1 U264 ( .B1(n532), .B2(n527), .A(n526), .ZN(n534) );
  INV_X1 U265 ( .A(n528), .ZN(n526) );
  NOR2_X1 U266 ( .A1(n518), .A2(n88), .ZN(n535) );
  INV_X1 U267 ( .A(n516), .ZN(n518) );
  OAI21_X1 U268 ( .B1(n517), .B2(n612), .A(n515), .ZN(n516) );
  AND2_X1 U269 ( .A1(n603), .A2(n569), .ZN(n600) );
  XNOR2_X1 U270 ( .A(n611), .B(n610), .ZN(n614) );
  NAND2_X1 U271 ( .A1(n608), .A2(n607), .ZN(n611) );
  INV_X1 U272 ( .A(n605), .ZN(n608) );
  NAND2_X1 U273 ( .A1(n416), .A2(n569), .ZN(n418) );
  INV_X1 U274 ( .A(n584), .ZN(n489) );
  AOI21_X1 U275 ( .B1(n536), .B2(n543), .A(n537), .ZN(n596) );
  NOR2_X1 U276 ( .A1(n603), .A2(n569), .ZN(n599) );
  NOR2_X1 U277 ( .A1(n463), .A2(n577), .ZN(n467) );
  NAND2_X1 U278 ( .A1(n463), .A2(n577), .ZN(n468) );
  AND2_X1 U279 ( .A1(n495), .A2(n326), .ZN(n500) );
  AOI21_X1 U280 ( .B1(n373), .B2(n86), .A(n372), .ZN(n377) );
  NOR2_X1 U281 ( .A1(n375), .A2(n374), .ZN(n376) );
  INV_X1 U282 ( .A(n418), .ZN(n414) );
  NOR2_X1 U283 ( .A1(n410), .A2(n567), .ZN(n405) );
  NOR2_X1 U284 ( .A1(n399), .A2(n577), .ZN(n403) );
  NAND2_X1 U285 ( .A1(n399), .A2(n577), .ZN(n402) );
  NAND2_X1 U286 ( .A1(n410), .A2(n567), .ZN(n406) );
  NOR2_X1 U287 ( .A1(n416), .A2(n569), .ZN(n419) );
  AOI211_X1 U288 ( .C1(n336), .C2(n372), .A(n335), .B(n374), .ZN(n337) );
  AOI21_X1 U289 ( .B1(n573), .B2(n572), .A(n571), .ZN(n622) );
  NOR2_X1 U290 ( .A1(n624), .A2(n326), .ZN(n625) );
  OAI21_X1 U291 ( .B1(n609), .B2(n605), .A(n512), .ZN(n514) );
  NOR2_X1 U292 ( .A1(n606), .A2(n511), .ZN(n512) );
  XNOR2_X1 U293 ( .A(n508), .B(n507), .ZN(n510) );
  OAI211_X1 U294 ( .C1(n503), .C2(n444), .A(n443), .B(n442), .ZN(n475) );
  INV_X1 U295 ( .A(n434), .ZN(n443) );
  OR2_X1 U296 ( .A1(n497), .A2(n435), .ZN(n444) );
  OR2_X1 U297 ( .A1(n426), .A2(n371), .ZN(n384) );
  INV_X1 U298 ( .A(n574), .ZN(n340) );
  NOR2_X1 U299 ( .A1(n330), .A2(n277), .ZN(n278) );
  INV_X1 U300 ( .A(n129), .ZN(n128) );
  AND2_X1 U301 ( .A1(n336), .A2(n86), .ZN(n83) );
  OR2_X1 U302 ( .A1(n423), .A2(n326), .ZN(n84) );
  AND2_X1 U303 ( .A1(n428), .A2(n381), .ZN(n85) );
  NAND2_X1 U304 ( .A1(n423), .A2(n326), .ZN(n420) );
  OR2_X1 U305 ( .A1(n368), .A2(n326), .ZN(n86) );
  INV_X1 U306 ( .A(n476), .ZN(n536) );
  NOR2_X1 U307 ( .A1(n540), .A2(n567), .ZN(n476) );
  OR2_X1 U308 ( .A1(n500), .A2(n498), .ZN(n87) );
  AND2_X1 U309 ( .A1(n517), .A2(n612), .ZN(n88) );
  OR2_X1 U310 ( .A1(n497), .A2(n498), .ZN(n89) );
  NOR2_X1 U311 ( .A1(n479), .A2(n567), .ZN(n481) );
  INV_X1 U312 ( .A(n481), .ZN(n413) );
  OR2_X1 U313 ( .A1(n568), .A2(n567), .ZN(n90) );
  OR2_X1 U314 ( .A1(n628), .A2(n627), .ZN(n91) );
  AND2_X1 U315 ( .A1(n565), .A2(n564), .ZN(n92) );
  INV_X1 U316 ( .A(n371), .ZN(n429) );
  NOR2_X1 U317 ( .A1(n432), .A2(n616), .ZN(n371) );
  OR2_X1 U318 ( .A1(n331), .A2(n330), .ZN(n93) );
  NOR2_X2 U319 ( .A1(reset), .A2(n666), .ZN(N4) );
  INV_X1 U320 ( .A(reset), .ZN(n639) );
  AND2_X1 U321 ( .A1(valid_in), .A2(n639), .ZN(N3) );
  AND2_X1 U322 ( .A1(enable_g), .A2(n639), .ZN(n685) );
  INV_X1 U323 ( .A(n616), .ZN(n132) );
  NOR2_X1 U324 ( .A1(enable_g), .A2(reset), .ZN(n630) );
  AOI22_X1 U325 ( .A1(n132), .A2(n685), .B1(n630), .B2(g[9]), .ZN(n94) );
  INV_X1 U326 ( .A(n94), .ZN(n54) );
  AOI21_X1 U327 ( .B1(enable_f), .B2(a_reg[0]), .A(reset), .ZN(n95) );
  INV_X1 U328 ( .A(n95), .ZN(n99) );
  NAND3_X1 U329 ( .A1(N4), .A2(a_reg[0]), .A3(n668), .ZN(n96) );
  OAI21_X1 U330 ( .B1(n668), .B2(n99), .A(n96), .ZN(n55) );
  OAI21_X1 U331 ( .B1(n667), .B2(f[1]), .A(f[0]), .ZN(n97) );
  OAI211_X1 U332 ( .C1(f[0]), .C2(f[1]), .A(N4), .B(n97), .ZN(n98) );
  OAI21_X1 U333 ( .B1(n664), .B2(n99), .A(n98), .ZN(n56) );
  NOR2_X1 U334 ( .A1(n673), .A2(n651), .ZN(n111) );
  AOI21_X1 U335 ( .B1(n673), .B2(n651), .A(n111), .ZN(n108) );
  NOR2_X1 U336 ( .A1(n667), .A2(n673), .ZN(n107) );
  NAND2_X1 U337 ( .A1(a_reg[0]), .A2(f[0]), .ZN(n100) );
  NOR2_X1 U338 ( .A1(n664), .A2(n100), .ZN(n106) );
  NAND2_X1 U339 ( .A1(n639), .A2(n666), .ZN(n285) );
  INV_X1 U340 ( .A(n285), .ZN(n295) );
  AOI22_X1 U341 ( .A1(n101), .A2(N4), .B1(f[2]), .B2(n295), .ZN(n679) );
  NAND2_X1 U342 ( .A1(n655), .A2(n129), .ZN(n102) );
  INV_X1 U343 ( .A(n326), .ZN(n184) );
  AOI22_X1 U344 ( .A1(n184), .A2(n685), .B1(n630), .B2(g[8]), .ZN(n104) );
  INV_X1 U345 ( .A(n104), .ZN(n53) );
  NAND2_X1 U346 ( .A1(a_reg[0]), .A2(a_reg[2]), .ZN(n105) );
  NAND3_X1 U347 ( .A1(f[3]), .A2(a_reg[0]), .A3(a_reg[2]), .ZN(n113) );
  INV_X1 U348 ( .A(n113), .ZN(n123) );
  AOI21_X1 U349 ( .B1(n669), .B2(n105), .A(n123), .ZN(n112) );
  FA_X1 U350 ( .A(n108), .B(n107), .CI(n106), .CO(n110), .S(n101) );
  AOI22_X1 U351 ( .A1(n109), .A2(N4), .B1(f[3]), .B2(n295), .ZN(n678) );
  NOR2_X1 U352 ( .A1(n674), .A2(n652), .ZN(n139) );
  AOI21_X1 U353 ( .B1(n674), .B2(n652), .A(n139), .ZN(n119) );
  NOR2_X1 U354 ( .A1(n667), .A2(n662), .ZN(n118) );
  NOR2_X1 U355 ( .A1(n674), .A2(n673), .ZN(n117) );
  FA_X1 U356 ( .A(n112), .B(n111), .CI(n110), .CO(n122), .S(n109) );
  INV_X1 U357 ( .A(n122), .ZN(n114) );
  NAND2_X1 U358 ( .A1(n113), .A2(n114), .ZN(n120) );
  OAI21_X1 U359 ( .B1(n114), .B2(n113), .A(n120), .ZN(n115) );
  XOR2_X1 U360 ( .A(n121), .B(n115), .Z(n116) );
  OAI22_X1 U361 ( .A1(n116), .A2(n294), .B1(n285), .B2(n652), .ZN(n59) );
  FA_X1 U362 ( .A(n119), .B(n118), .CI(n117), .CO(n135), .S(n121) );
  AOI22_X1 U363 ( .A1(n123), .A2(n122), .B1(n121), .B2(n120), .ZN(n124) );
  INV_X1 U364 ( .A(n124), .ZN(n136) );
  XOR2_X1 U365 ( .A(n135), .B(n136), .Z(n126) );
  NAND2_X1 U366 ( .A1(a_reg[1]), .A2(a_reg[3]), .ZN(n125) );
  NOR3_X1 U367 ( .A1(n663), .A2(n673), .A3(n662), .ZN(n147) );
  AOI21_X1 U368 ( .B1(n663), .B2(n125), .A(n147), .ZN(n140) );
  NOR2_X1 U369 ( .A1(n667), .A2(n661), .ZN(n138) );
  XNOR2_X1 U370 ( .A(n126), .B(n134), .ZN(n127) );
  OAI22_X1 U371 ( .A1(n127), .A2(n294), .B1(n285), .B2(n663), .ZN(n60) );
  AOI222_X1 U372 ( .A1(f[17]), .A2(n326), .B1(f[17]), .B2(f[16]), .C1(n129), 
        .C2(n184), .ZN(n190) );
  NOR2_X1 U373 ( .A1(f[15]), .A2(f[14]), .ZN(n185) );
  INV_X1 U374 ( .A(n185), .ZN(n186) );
  AOI22_X1 U375 ( .A1(f[16]), .A2(n326), .B1(n186), .B2(n656), .ZN(n191) );
  AND2_X1 U376 ( .A1(n132), .A2(n190), .ZN(n131) );
  OAI221_X1 U377 ( .B1(f[18]), .B2(n129), .C1(n655), .C2(n128), .A(f[19]), 
        .ZN(n130) );
  OAI221_X1 U378 ( .B1(n132), .B2(n190), .C1(n191), .C2(n131), .A(n130), .ZN(
        n257) );
  AOI22_X1 U379 ( .A1(n257), .A2(n685), .B1(n630), .B2(g[7]), .ZN(n133) );
  INV_X1 U380 ( .A(n133), .ZN(n52) );
  NOR2_X1 U381 ( .A1(n661), .A2(n673), .ZN(n144) );
  NOR2_X1 U382 ( .A1(n667), .A2(n672), .ZN(n143) );
  NOR2_X1 U383 ( .A1(n674), .A2(n662), .ZN(n142) );
  NOR2_X1 U384 ( .A1(n662), .A2(n653), .ZN(n161) );
  AOI21_X1 U385 ( .B1(n662), .B2(n653), .A(n161), .ZN(n146) );
  OAI222_X1 U386 ( .A1(n136), .A2(n135), .B1(n136), .B2(n134), .C1(n135), .C2(
        n134), .ZN(n137) );
  INV_X1 U387 ( .A(n137), .ZN(n150) );
  FA_X1 U388 ( .A(n140), .B(n139), .CI(n138), .CO(n149), .S(n134) );
  AOI22_X1 U389 ( .A1(n141), .A2(N4), .B1(f[6]), .B2(n295), .ZN(n677) );
  NOR2_X1 U390 ( .A1(n667), .A2(n659), .ZN(n160) );
  NOR2_X1 U391 ( .A1(n673), .A2(n672), .ZN(n159) );
  FA_X1 U392 ( .A(n144), .B(n143), .CI(n142), .CO(n157), .S(n148) );
  NAND2_X1 U393 ( .A1(a_reg[2]), .A2(a_reg[4]), .ZN(n145) );
  NOR3_X1 U394 ( .A1(n674), .A2(n665), .A3(n661), .ZN(n168) );
  AOI21_X1 U395 ( .B1(n665), .B2(n145), .A(n168), .ZN(n156) );
  FA_X1 U396 ( .A(n148), .B(n147), .CI(n146), .CO(n154), .S(n151) );
  FA_X1 U397 ( .A(n151), .B(n150), .CI(n149), .CO(n153), .S(n141) );
  AOI22_X1 U398 ( .A1(n152), .A2(N4), .B1(f[7]), .B2(n295), .ZN(n676) );
  FA_X1 U399 ( .A(n155), .B(n154), .CI(n153), .CO(n171), .S(n152) );
  FA_X1 U400 ( .A(n158), .B(n157), .CI(n156), .CO(n172), .S(n155) );
  NOR2_X1 U401 ( .A1(n172), .A2(n171), .ZN(n175) );
  AOI21_X1 U402 ( .B1(n171), .B2(n172), .A(n175), .ZN(n163) );
  NOR2_X1 U403 ( .A1(n654), .A2(n661), .ZN(n206) );
  AOI21_X1 U404 ( .B1(n654), .B2(n661), .A(n206), .ZN(n170) );
  NOR2_X1 U405 ( .A1(n661), .A2(n662), .ZN(n169) );
  NOR2_X1 U406 ( .A1(n674), .A2(n672), .ZN(n167) );
  NOR2_X1 U407 ( .A1(n667), .A2(n660), .ZN(n166) );
  NOR2_X1 U408 ( .A1(n659), .A2(n673), .ZN(n165) );
  FA_X1 U409 ( .A(n161), .B(n160), .CI(n159), .CO(n176), .S(n158) );
  INV_X1 U410 ( .A(n162), .ZN(n174) );
  XOR2_X1 U411 ( .A(n163), .B(n174), .Z(n164) );
  OAI22_X1 U412 ( .A1(n164), .A2(n294), .B1(n285), .B2(n654), .ZN(n63) );
  NOR2_X1 U413 ( .A1(n660), .A2(n673), .ZN(n205) );
  FA_X1 U414 ( .A(n167), .B(n166), .CI(n165), .CO(n204), .S(n177) );
  FA_X1 U415 ( .A(n170), .B(n169), .CI(n168), .CO(n199), .S(n178) );
  NOR2_X1 U416 ( .A1(n674), .A2(n659), .ZN(n202) );
  NOR2_X1 U417 ( .A1(n662), .A2(n672), .ZN(n201) );
  NAND2_X1 U418 ( .A1(n172), .A2(n171), .ZN(n173) );
  OAI21_X1 U419 ( .B1(n175), .B2(n174), .A(n173), .ZN(n196) );
  FA_X1 U420 ( .A(n178), .B(n177), .CI(n176), .CO(n195), .S(n162) );
  AOI22_X1 U421 ( .A1(n179), .A2(N4), .B1(f[9]), .B2(n295), .ZN(n180) );
  INV_X1 U422 ( .A(n180), .ZN(n64) );
  NAND2_X1 U423 ( .A1(n267), .A2(n184), .ZN(n263) );
  INV_X1 U424 ( .A(n263), .ZN(n183) );
  NOR2_X1 U425 ( .A1(f[12]), .A2(f[13]), .ZN(n258) );
  INV_X1 U426 ( .A(n258), .ZN(n259) );
  AOI22_X1 U427 ( .A1(f[14]), .A2(n569), .B1(n259), .B2(n658), .ZN(n265) );
  NAND2_X1 U428 ( .A1(n326), .A2(n182), .ZN(n262) );
  OAI21_X1 U429 ( .B1(n183), .B2(n265), .A(n262), .ZN(n273) );
  AOI22_X1 U430 ( .A1(f[16]), .A2(n326), .B1(n184), .B2(n656), .ZN(n188) );
  AOI22_X1 U431 ( .A1(f[16]), .A2(n186), .B1(n185), .B2(n656), .ZN(n187) );
  AOI22_X1 U432 ( .A1(n569), .A2(n188), .B1(n187), .B2(n257), .ZN(n276) );
  OR2_X1 U433 ( .A1(n616), .A2(n276), .ZN(n193) );
  AOI21_X1 U434 ( .B1(n257), .B2(n190), .A(n191), .ZN(n189) );
  AOI211_X1 U435 ( .C1(n191), .C2(n190), .A(n189), .B(n616), .ZN(n192) );
  AOI221_X4 U436 ( .B1(n273), .B2(n193), .C1(n616), .C2(n276), .A(n192), .ZN(
        n567) );
  AOI22_X1 U437 ( .A1(n253), .A2(n685), .B1(n630), .B2(g[6]), .ZN(n194) );
  INV_X1 U438 ( .A(n194), .ZN(n51) );
  FA_X1 U439 ( .A(n197), .B(n196), .CI(n195), .CO(n213), .S(n179) );
  FA_X1 U440 ( .A(n200), .B(n199), .CI(n198), .CO(n214), .S(n197) );
  NOR2_X1 U441 ( .A1(n214), .A2(n213), .ZN(n217) );
  AOI21_X1 U442 ( .B1(n213), .B2(n214), .A(n217), .ZN(n208) );
  NOR2_X1 U443 ( .A1(n674), .A2(n660), .ZN(n212) );
  NOR2_X1 U444 ( .A1(n659), .A2(n662), .ZN(n211) );
  FA_X1 U445 ( .A(f[9]), .B(n202), .CI(n201), .CO(n210), .S(n198) );
  NAND2_X1 U446 ( .A1(n661), .A2(a_reg[5]), .ZN(n203) );
  XOR2_X1 U447 ( .A(n203), .B(n650), .Z(n219) );
  FA_X1 U448 ( .A(n206), .B(n205), .CI(n204), .CO(n218), .S(n200) );
  INV_X1 U449 ( .A(n207), .ZN(n216) );
  XOR2_X1 U450 ( .A(n208), .B(n216), .Z(n209) );
  OAI22_X1 U451 ( .A1(n209), .A2(n294), .B1(n285), .B2(n650), .ZN(n65) );
  NOR2_X1 U452 ( .A1(n660), .A2(n662), .ZN(n225) );
  NOR2_X1 U453 ( .A1(n659), .A2(n661), .ZN(n224) );
  AOI21_X1 U454 ( .B1(n650), .B2(n661), .A(n672), .ZN(n227) );
  FA_X1 U455 ( .A(n212), .B(n211), .CI(n210), .CO(n226), .S(n220) );
  NAND2_X1 U456 ( .A1(n214), .A2(n213), .ZN(n215) );
  OAI21_X1 U457 ( .B1(n217), .B2(n216), .A(n215), .ZN(n230) );
  FA_X1 U458 ( .A(n220), .B(n219), .CI(n218), .CO(n229), .S(n207) );
  AOI22_X1 U459 ( .A1(n221), .A2(N4), .B1(f[11]), .B2(n295), .ZN(n222) );
  INV_X1 U460 ( .A(n222), .ZN(n66) );
  NOR2_X1 U461 ( .A1(a_reg[5]), .A2(n659), .ZN(n223) );
  XOR2_X1 U462 ( .A(f[12]), .B(n223), .Z(n235) );
  NOR2_X1 U463 ( .A1(n660), .A2(n661), .ZN(n234) );
  FA_X1 U464 ( .A(f[11]), .B(n225), .CI(n224), .CO(n233), .S(n228) );
  FA_X1 U465 ( .A(n228), .B(n227), .CI(n226), .CO(n237), .S(n231) );
  FA_X1 U466 ( .A(n231), .B(n230), .CI(n229), .CO(n236), .S(n221) );
  AOI22_X1 U467 ( .A1(n232), .A2(N4), .B1(f[12]), .B2(n295), .ZN(n675) );
  AOI21_X1 U468 ( .B1(n672), .B2(n657), .A(n659), .ZN(n243) );
  NOR2_X1 U469 ( .A1(n660), .A2(n672), .ZN(n242) );
  FA_X1 U470 ( .A(n235), .B(n234), .CI(n233), .CO(n247), .S(n238) );
  FA_X1 U471 ( .A(n238), .B(n237), .CI(n236), .CO(n246), .S(n232) );
  NAND2_X1 U472 ( .A1(n247), .A2(n246), .ZN(n239) );
  OR2_X1 U473 ( .A1(n247), .A2(n246), .ZN(n244) );
  NAND2_X1 U474 ( .A1(n239), .A2(n244), .ZN(n240) );
  XOR2_X1 U475 ( .A(n245), .B(n240), .Z(n241) );
  OAI22_X1 U476 ( .A1(n241), .A2(n294), .B1(n285), .B2(n670), .ZN(n68) );
  FA_X1 U477 ( .A(f[13]), .B(n243), .CI(n242), .CO(n283), .S(n245) );
  AOI22_X1 U478 ( .A1(n247), .A2(n246), .B1(n245), .B2(n244), .ZN(n248) );
  INV_X1 U479 ( .A(n248), .ZN(n281) );
  XOR2_X1 U480 ( .A(n283), .B(n281), .Z(n250) );
  NAND2_X1 U481 ( .A1(a_reg[7]), .A2(n659), .ZN(n249) );
  XOR2_X1 U482 ( .A(n658), .B(n249), .Z(n282) );
  XNOR2_X1 U483 ( .A(n250), .B(n282), .ZN(n251) );
  OAI22_X1 U484 ( .A1(n251), .A2(n294), .B1(n285), .B2(n658), .ZN(n69) );
  NAND2_X1 U485 ( .A1(n567), .A2(n657), .ZN(n252) );
  OAI21_X1 U486 ( .B1(n567), .B2(n657), .A(n252), .ZN(n254) );
  INV_X1 U487 ( .A(n567), .ZN(n253) );
  NAND2_X1 U488 ( .A1(n254), .A2(n253), .ZN(n304) );
  OR2_X1 U489 ( .A1(f[10]), .A2(f[11]), .ZN(n306) );
  NAND2_X1 U490 ( .A1(n304), .A2(n306), .ZN(n255) );
  NAND2_X1 U491 ( .A1(n307), .A2(n567), .ZN(n303) );
  INV_X1 U492 ( .A(n329), .ZN(n271) );
  OAI21_X1 U493 ( .B1(n567), .B2(f[12]), .A(f[13]), .ZN(n256) );
  OAI21_X1 U494 ( .B1(n567), .B2(n259), .A(n256), .ZN(n324) );
  AOI22_X1 U495 ( .A1(f[14]), .A2(n569), .B1(n257), .B2(n658), .ZN(n261) );
  AOI22_X1 U496 ( .A1(f[14]), .A2(n259), .B1(n258), .B2(n658), .ZN(n260) );
  AOI22_X1 U497 ( .A1(n567), .A2(n261), .B1(n260), .B2(n253), .ZN(n319) );
  INV_X1 U498 ( .A(n327), .ZN(n270) );
  NAND2_X1 U499 ( .A1(n263), .A2(n262), .ZN(n264) );
  XNOR2_X1 U500 ( .A(n265), .B(n264), .ZN(n266) );
  AOI22_X1 U501 ( .A1(n567), .A2(n267), .B1(n266), .B2(n253), .ZN(n333) );
  NAND2_X1 U502 ( .A1(n327), .A2(n328), .ZN(n268) );
  OAI211_X1 U503 ( .C1(n271), .C2(n270), .A(n269), .B(n268), .ZN(n279) );
  NAND2_X1 U504 ( .A1(n616), .A2(n273), .ZN(n272) );
  OAI211_X1 U505 ( .C1(n273), .C2(n616), .A(n272), .B(n253), .ZN(n275) );
  NAND2_X1 U506 ( .A1(n275), .A2(n276), .ZN(n274) );
  OAI21_X1 U507 ( .B1(n276), .B2(n275), .A(n274), .ZN(n277) );
  NAND2_X1 U508 ( .A1(n279), .A2(n278), .ZN(n300) );
  AOI22_X1 U509 ( .A1(n300), .A2(n685), .B1(n630), .B2(g[5]), .ZN(n280) );
  INV_X1 U510 ( .A(n280), .ZN(n50) );
  AOI222_X1 U511 ( .A1(n283), .A2(n282), .B1(n283), .B2(n281), .C1(n282), .C2(
        n281), .ZN(n287) );
  OAI21_X1 U512 ( .B1(f[14]), .B2(a_reg[6]), .A(a_reg[7]), .ZN(n288) );
  XOR2_X1 U513 ( .A(f[15]), .B(n288), .Z(n284) );
  XNOR2_X1 U514 ( .A(n287), .B(n284), .ZN(n286) );
  OAI22_X1 U515 ( .A1(n286), .A2(n294), .B1(n285), .B2(n648), .ZN(n70) );
  INV_X1 U516 ( .A(n288), .ZN(n290) );
  OAI21_X1 U517 ( .B1(n288), .B2(n648), .A(n287), .ZN(n289) );
  OAI21_X1 U518 ( .B1(f[15]), .B2(n290), .A(n289), .ZN(n293) );
  OAI21_X1 U519 ( .B1(n293), .B2(n666), .A(n639), .ZN(n292) );
  NOR2_X1 U520 ( .A1(n294), .A2(n293), .ZN(n297) );
  NAND2_X1 U521 ( .A1(n656), .A2(n297), .ZN(n291) );
  OAI21_X1 U522 ( .B1(n292), .B2(n656), .A(n291), .ZN(n71) );
  INV_X1 U523 ( .A(n293), .ZN(n634) );
  AOI21_X1 U524 ( .B1(n634), .B2(f[16]), .A(n294), .ZN(n296) );
  OAI21_X1 U525 ( .B1(n296), .B2(n295), .A(f[17]), .ZN(n299) );
  NAND3_X1 U526 ( .A1(n671), .A2(f[16]), .A3(n297), .ZN(n298) );
  NAND2_X1 U527 ( .A1(n299), .A2(n298), .ZN(n72) );
  AOI22_X1 U528 ( .A1(n300), .A2(f[10]), .B1(n650), .B2(n577), .ZN(n347) );
  OR2_X1 U529 ( .A1(f[8]), .A2(f[9]), .ZN(n346) );
  OAI21_X1 U530 ( .B1(n577), .B2(f[10]), .A(f[11]), .ZN(n302) );
  OAI21_X1 U531 ( .B1(n577), .B2(n306), .A(n302), .ZN(n363) );
  NAND2_X1 U532 ( .A1(n304), .A2(n303), .ZN(n305) );
  MUX2_X1 U533 ( .A(n308), .B(n307), .S(n577), .Z(n357) );
  MUX2_X1 U534 ( .A(n320), .B(n319), .S(n577), .Z(n378) );
  XNOR2_X1 U535 ( .A(n323), .B(n329), .ZN(n325) );
  MUX2_X1 U536 ( .A(n325), .B(n324), .S(n577), .Z(n368) );
  XNOR2_X1 U537 ( .A(n332), .B(n93), .ZN(n334) );
  MUX2_X1 U538 ( .A(n334), .B(n333), .S(n577), .Z(n335) );
  INV_X1 U539 ( .A(n337), .ZN(n338) );
  AOI22_X1 U540 ( .A1(n340), .A2(n685), .B1(n630), .B2(g[4]), .ZN(n339) );
  INV_X1 U541 ( .A(n339), .ZN(n49) );
  AOI22_X1 U542 ( .A1(n340), .A2(f[8]), .B1(n654), .B2(n574), .ZN(n391) );
  OR2_X1 U543 ( .A1(f[6]), .A2(f[7]), .ZN(n390) );
  OAI21_X1 U544 ( .B1(n574), .B2(f[8]), .A(f[9]), .ZN(n342) );
  OAI21_X1 U545 ( .B1(n574), .B2(n346), .A(n342), .ZN(n399) );
  NAND2_X1 U546 ( .A1(n344), .A2(n343), .ZN(n345) );
  MUX2_X1 U547 ( .A(n348), .B(n347), .S(n574), .Z(n410) );
  MUX2_X1 U548 ( .A(n358), .B(n357), .S(n574), .Z(n423) );
  XNOR2_X1 U549 ( .A(n362), .B(n361), .ZN(n364) );
  XNOR2_X1 U550 ( .A(n373), .B(n367), .ZN(n369) );
  MUX2_X1 U551 ( .A(n369), .B(n368), .S(n574), .Z(n432) );
  NAND2_X1 U552 ( .A1(n414), .A2(n84), .ZN(n370) );
  AND2_X1 U553 ( .A1(n370), .A2(n420), .ZN(n425) );
  MUX2_X1 U554 ( .A(n379), .B(n378), .S(n574), .Z(n380) );
  OAI21_X1 U555 ( .B1(n425), .B2(n371), .A(n85), .ZN(n382) );
  INV_X1 U556 ( .A(n382), .ZN(n383) );
  OAI21_X1 U557 ( .B1(n427), .B2(n384), .A(n383), .ZN(n393) );
  AOI22_X1 U558 ( .A1(n393), .A2(n685), .B1(n630), .B2(g[3]), .ZN(n385) );
  INV_X1 U559 ( .A(n385), .ZN(n48) );
  OAI21_X1 U560 ( .B1(n529), .B2(f[6]), .A(f[7]), .ZN(n386) );
  OAI21_X1 U561 ( .B1(n529), .B2(n390), .A(n386), .ZN(n460) );
  NAND2_X1 U562 ( .A1(n388), .A2(n387), .ZN(n389) );
  MUX2_X1 U563 ( .A(n392), .B(n391), .S(n529), .Z(n463) );
  NOR2_X1 U564 ( .A1(n465), .A2(n467), .ZN(n396) );
  AOI22_X1 U565 ( .A1(n393), .A2(f[6]), .B1(n653), .B2(n529), .ZN(n451) );
  OR2_X1 U566 ( .A1(f[4]), .A2(f[5]), .ZN(n450) );
  INV_X1 U567 ( .A(n403), .ZN(n397) );
  NAND2_X1 U568 ( .A1(n397), .A2(n402), .ZN(n398) );
  MUX2_X1 U569 ( .A(n400), .B(n399), .S(n529), .Z(n479) );
  MUX2_X1 U570 ( .A(n411), .B(n410), .S(n529), .Z(n487) );
  NAND2_X1 U571 ( .A1(n412), .A2(n257), .ZN(n484) );
  XNOR2_X1 U572 ( .A(n427), .B(n415), .ZN(n417) );
  MUX2_X1 U573 ( .A(n417), .B(n416), .S(n529), .Z(n495) );
  OAI21_X1 U574 ( .B1(n427), .B2(n419), .A(n418), .ZN(n422) );
  NAND2_X1 U575 ( .A1(n84), .A2(n420), .ZN(n421) );
  MUX2_X1 U576 ( .A(n424), .B(n423), .S(n529), .Z(n509) );
  OAI21_X1 U577 ( .B1(n427), .B2(n426), .A(n425), .ZN(n431) );
  MUX2_X1 U578 ( .A(n433), .B(n432), .S(n529), .Z(n434) );
  INV_X1 U579 ( .A(n482), .ZN(n437) );
  INV_X1 U580 ( .A(n483), .ZN(n436) );
  AOI21_X1 U581 ( .B1(n484), .B2(n437), .A(n436), .ZN(n499) );
  INV_X1 U582 ( .A(n499), .ZN(n440) );
  AOI21_X1 U583 ( .B1(n441), .B2(n440), .A(n439), .ZN(n442) );
  AOI22_X1 U584 ( .A1(n475), .A2(n685), .B1(n630), .B2(g[2]), .ZN(n445) );
  INV_X1 U585 ( .A(n445), .ZN(n47) );
  OAI21_X1 U586 ( .B1(n527), .B2(f[4]), .A(f[5]), .ZN(n446) );
  OAI21_X1 U587 ( .B1(n527), .B2(n450), .A(n446), .ZN(n561) );
  NAND2_X1 U588 ( .A1(n448), .A2(n447), .ZN(n449) );
  MUX2_X1 U589 ( .A(n452), .B(n451), .S(n527), .Z(n555) );
  AOI22_X1 U590 ( .A1(n475), .A2(f[4]), .B1(n652), .B2(n527), .ZN(n524) );
  OR2_X1 U591 ( .A1(f[2]), .A2(f[3]), .ZN(n523) );
  NAND2_X1 U592 ( .A1(n524), .A2(n527), .ZN(n520) );
  AOI21_X1 U593 ( .B1(n558), .B2(n552), .A(n550), .ZN(n455) );
  MUX2_X1 U594 ( .A(n461), .B(n460), .S(n527), .Z(n547) );
  INV_X1 U595 ( .A(n547), .ZN(n462) );
  INV_X1 U596 ( .A(n467), .ZN(n469) );
  NAND2_X1 U597 ( .A1(n544), .A2(n536), .ZN(n595) );
  NAND2_X1 U598 ( .A1(n413), .A2(n482), .ZN(n478) );
  MUX2_X1 U599 ( .A(n480), .B(n479), .S(n527), .Z(n603) );
  MUX2_X1 U600 ( .A(n488), .B(n487), .S(n527), .Z(n593) );
  AOI21_X1 U601 ( .B1(n600), .B2(n584), .A(n583), .ZN(n490) );
  OAI21_X1 U602 ( .B1(n503), .B2(n497), .A(n499), .ZN(n494) );
  MUX2_X1 U603 ( .A(n496), .B(n495), .S(n527), .Z(n613) );
  NOR2_X1 U604 ( .A1(n499), .A2(n498), .ZN(n501) );
  INV_X1 U605 ( .A(n504), .ZN(n506) );
  MUX2_X1 U606 ( .A(n510), .B(n509), .S(n527), .Z(n511) );
  AOI22_X1 U607 ( .A1(n514), .A2(n685), .B1(n630), .B2(g[1]), .ZN(n513) );
  INV_X1 U608 ( .A(n513), .ZN(n46) );
  AOI22_X1 U609 ( .A1(n514), .A2(f[2]), .B1(n651), .B2(n612), .ZN(n517) );
  OR2_X1 U610 ( .A1(f[0]), .A2(f[1]), .ZN(n515) );
  OAI21_X1 U611 ( .B1(n612), .B2(f[2]), .A(f[3]), .ZN(n519) );
  OAI21_X1 U612 ( .B1(n612), .B2(n523), .A(n519), .ZN(n532) );
  MUX2_X1 U613 ( .A(n525), .B(n524), .S(n612), .Z(n530) );
  OAI21_X1 U614 ( .B1(n535), .B2(n534), .A(n533), .ZN(n566) );
  MUX2_X1 U615 ( .A(n541), .B(n540), .S(n612), .Z(n570) );
  INV_X1 U616 ( .A(n570), .ZN(n542) );
  INV_X1 U617 ( .A(n543), .ZN(n545) );
  NAND2_X1 U618 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U619 ( .A(n598), .B(n546), .ZN(n548) );
  MUX2_X1 U620 ( .A(n548), .B(n547), .S(n612), .Z(n568) );
  INV_X1 U621 ( .A(n581), .ZN(n565) );
  INV_X1 U622 ( .A(n558), .ZN(n549) );
  INV_X1 U623 ( .A(n550), .ZN(n551) );
  MUX2_X1 U624 ( .A(n556), .B(n555), .S(n612), .Z(n578) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n562) );
  MUX2_X1 U627 ( .A(n562), .B(n561), .S(n612), .Z(n575) );
  NAND2_X1 U628 ( .A1(n566), .A2(n92), .ZN(n623) );
  OR2_X1 U629 ( .A1(n582), .A2(n581), .ZN(n621) );
  INV_X1 U630 ( .A(n583), .ZN(n585) );
  INV_X1 U631 ( .A(n599), .ZN(n587) );
  INV_X1 U632 ( .A(n595), .ZN(n586) );
  NAND3_X1 U633 ( .A1(n587), .A2(n586), .A3(n598), .ZN(n590) );
  NOR2_X1 U634 ( .A1(n596), .A2(n599), .ZN(n588) );
  MUX2_X1 U635 ( .A(n594), .B(n593), .S(n612), .Z(n617) );
  INV_X1 U636 ( .A(n596), .ZN(n597) );
  MUX2_X1 U637 ( .A(n604), .B(n603), .S(n612), .Z(n624) );
  INV_X1 U638 ( .A(n609), .ZN(n610) );
  MUX2_X1 U639 ( .A(n614), .B(n613), .S(n612), .Z(n615) );
  INV_X1 U640 ( .A(n628), .ZN(n620) );
  NAND4_X1 U641 ( .A1(n623), .A2(n622), .A3(n621), .A4(n620), .ZN(n629) );
  NOR2_X1 U642 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U643 ( .A1(n629), .A2(n91), .ZN(n633) );
  INV_X1 U644 ( .A(n685), .ZN(n632) );
  NAND2_X1 U645 ( .A1(n630), .A2(g[0]), .ZN(n631) );
  OAI21_X1 U646 ( .B1(n633), .B2(n632), .A(n631), .ZN(n45) );
  NAND3_X1 U647 ( .A1(n634), .A2(f[17]), .A3(f[16]), .ZN(n636) );
  OAI21_X1 U648 ( .B1(n636), .B2(f[19]), .A(f[18]), .ZN(n635) );
  OAI211_X1 U649 ( .C1(f[18]), .C2(f[19]), .A(n635), .B(N4), .ZN(n638) );
  INV_X1 U650 ( .A(n636), .ZN(n641) );
  NAND2_X1 U651 ( .A1(n641), .A2(enable_f), .ZN(n640) );
  NAND3_X1 U652 ( .A1(n640), .A2(f[19]), .A3(n639), .ZN(n637) );
  NAND2_X1 U653 ( .A1(n638), .A2(n637), .ZN(n74) );
  NAND3_X1 U654 ( .A1(n640), .A2(f[18]), .A3(n639), .ZN(n643) );
  NAND3_X1 U655 ( .A1(n641), .A2(N4), .A3(n655), .ZN(n642) );
  NAND2_X1 U656 ( .A1(n643), .A2(n642), .ZN(n73) );
  NOR2_X1 U657 ( .A1(reset), .A2(valid_in), .ZN(n647) );
  AOI22_X1 U658 ( .A1(a_reg[7]), .A2(n647), .B1(N3), .B2(a[7]), .ZN(n680) );
  AOI22_X1 U659 ( .A1(a_reg[6]), .A2(n647), .B1(N3), .B2(a[6]), .ZN(n681) );
  AOI22_X1 U660 ( .A1(n647), .A2(a_reg[5]), .B1(N3), .B2(a[5]), .ZN(n644) );
  INV_X1 U661 ( .A(n644), .ZN(n80) );
  AOI22_X1 U662 ( .A1(a_reg[4]), .A2(n647), .B1(N3), .B2(a[4]), .ZN(n682) );
  AOI22_X1 U663 ( .A1(a_reg[3]), .A2(n647), .B1(N3), .B2(a[3]), .ZN(n683) );
  AOI22_X1 U664 ( .A1(a_reg[2]), .A2(n647), .B1(N3), .B2(a[2]), .ZN(n645) );
  INV_X1 U665 ( .A(n645), .ZN(n77) );
  AOI22_X1 U666 ( .A1(a_reg[1]), .A2(n647), .B1(N3), .B2(a[1]), .ZN(n646) );
  INV_X1 U667 ( .A(n646), .ZN(n76) );
  AOI22_X1 U668 ( .A1(a_reg[0]), .A2(n647), .B1(N3), .B2(a[0]), .ZN(n684) );
endmodule

